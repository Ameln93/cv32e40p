// Copyright 2018 Robert Balas <balasr@student.ethz.ch>
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Wrapper for a RI5CY testbench, containing RI5CY, Memory and stdout peripheral
// Contributor: Robert Balas <balasr@student.ethz.ch>

module riscv_wrapper
#(parameter INSTR_RDATA_WIDTH = 128,
  parameter RAM_ADDR_WIDTH    = 20,
  parameter BOOT_ADDR         = 'h80,
  parameter PULP_SECURE       = 1,
  parameter VPU               = 1,
  parameter VLEN              = 128,
  parameter LANES             = 2
)(
  input logic         clk_i,
  input logic         rst_ni,

  input logic         fetch_enable_i,
  output logic        tests_passed_o,
  output logic        tests_failed_o,
  output logic [31:0] exit_value_o,
  output logic        exit_valid_o
);

// signals connecting core to memory
logic                         instr_req;
logic                         instr_gnt;
logic                         instr_rvalid;
logic [31:0]                  instr_addr;
logic [INSTR_RDATA_WIDTH-1:0] instr_rdata;

logic                         apu_req;
logic                         apu_gnt;
logic [2:0][31:0]             apu_operands;
logic                         apu_rvalid;
logic [31:0]                  apu_rdata;



logic                         data_cpu_req;
logic                         data_cpu_gnt;
logic                         data_cpu_rvalid;
logic [31:0]                  data_cpu_addr;
logic                         data_cpu_we;
logic [3:0]                   data_cpu_be;
logic [31:0]                  data_cpu_rdata;
logic [31:0]                  data_cpu_wdata;

logic                         data_vpu_req;
logic                         data_vpu_gnt;
logic                         data_vpu_rvalid;
logic [31:0]                  data_vpu_addr;
logic                         data_vpu_we;
logic [3:0]                   data_vpu_be;
logic [31:0]                  data_vpu_rdata;
logic [31:0]                  data_vpu_wdata;


logic                         data_gnt;
logic [31:0]                  data_rdata;
logic                         data_rvalid;
logic                         data_req;
logic [31:0]                  data_addr;
logic                         data_we;
logic [3:0]                   data_be;
logic [31:0]                  data_wdata;


// signals to debug unit
logic                         debug_req_i;

// irq signals (not used)
logic                         irq;
logic [0:4]                   irq_id_in;
logic                         irq_ack;
logic [0:4]                   irq_id_out;
logic                         irq_sec;


// interrupts (only timer for now)
assign irq_sec     = '0;

assign debug_req_i = 1'b0;

// instantiate the core
riscv_core
#(.INSTR_RDATA_WIDTH (INSTR_RDATA_WIDTH),
  .PULP_SECURE(PULP_SECURE),
  .VPU(1),
  .VLEN(VLEN),
  .FPU(0)
)
riscv_core_i
(
  .clk_i                  ( clk_i                 ),
  .rst_ni                 ( rst_ni                ),

  .clock_en_i             ( '1                    ),
  .test_en_i              ( '0                    ),

  .boot_addr_i            ( BOOT_ADDR             ),
  .core_id_i              ( 4'h0                  ),
  .cluster_id_i           ( 6'h0                  ),

  .instr_addr_o           ( instr_addr            ),
  .instr_req_o            ( instr_req             ),
  .instr_rdata_i          ( instr_rdata           ),
  .instr_gnt_i            ( instr_gnt             ),
  .instr_rvalid_i         ( instr_rvalid          ),

  .data_addr_o            ( data_cpu_addr         ),
  .data_wdata_o           ( data_cpu_wdata        ),
  .data_we_o              ( data_cpu_we           ),
  .data_req_o             ( data_cpu_req          ),
  .data_be_o              ( data_cpu_be           ),
  .data_rdata_i           ( data_cpu_rdata        ),
  .data_gnt_i             ( data_cpu_gnt          ),
  .data_rvalid_i          ( data_cpu_rvalid       ),

  .apu_master_req_o       ( apu_req               ),
  .apu_master_ready_o     (/*cpu is always ready*/),
  .apu_master_gnt_i       ( apu_gnt               ),
  .apu_master_operands_o  ( apu_operands          ),
  .apu_master_op_o        (/*not used by vpu*/    ),
  .apu_master_type_o      (/*not used by vpu*/    ),
  .apu_master_flags_o     (/*not used by vpu*/    ),
  .apu_master_valid_i     ( apu_rvalid            ),
  .apu_master_result_i    ( apu_rcsr              ),
  .apu_master_flags_i     ( /*not used by vpu*/   ),

  .irq_i                  ( irq                   ),
  .irq_id_i               ( irq_id_in             ),
  .irq_ack_o              ( irq_ack               ),
  .irq_id_o               ( irq_id_out            ),
  .irq_sec_i              ( irq_sec               ),

  .sec_lvl_o              ( sec_lvl_o             ),

  .debug_req_i            ( debug_req_i           ),

  .fetch_enable_i         ( fetch_enable_i        ),
  .core_busy_o            ( core_busy_o           ),

  .ext_perf_counters_i    (                       ),
  .fregfile_disable_i     ( 1'b0                  )
);

vpu_core #(
  .VLEN   (VLEN),
  .LANES  (LANES),
  .ELEN   (32)
)
vpu_i
(
  .clk_i                  ( clk_i                   ),
  .rst_ni                 ( rst_ni                  ),

  // insn interface
  .insn_req_i             ( apu_req                 ),
  .insn_gnt_o             ( apu_gnt                 ),
  .insn_data_i            ( apu_operands[0]         ),
  .insn_csr_i             ( apu_operands[1]         ),
  .insn_addr_i            ( apu_operands[2]         ),
  .insn_rvalid_o          ( apu_rvalid              ),
  .insn_rcsr_o            ( apu_rcsr                ),

  // data interface
  .data_req_o             ( data_vpu_req            ),
  .data_addr_o            ( data_vpu_addr           ),
  .data_be_o              ( data_vpu_be             ),
  .data_we_o              ( data_vpu_we             ),
  .data_wdata_o           ( data_vpu_wdata          ),
  .data_gnt_i             ( data_vpu_gnt            ),
  .data_rvalid_i          ( data_vpu_rvalid         ),
  .data_rdata_i           ( data_vpu_rdata          ),

  .dbg_ex_wb_hs_o         (                         ),
  .dbg_ex_wb_en_o         (                         ),
  .dbg_if_id_en_o         (                         ),
  .dbg_alu_carry_o        (                         ),
  .dbg_arith_result_o     (                         ),
  .dbg_arith_valid_o      (                         ),
  .dbg_byte_enable_o      (                         ),
  .dbg_iteration_o        (                         ),
  .dbg_insn_complete_o    (                         )
);

obi_arbiter arbiter_i
(
  .clk_i                  ( clk_i                  ),
  .rst_ni                 ( rst_ni                 ),
  // input slave a vpu (priorized
  .s_req_a_i              ( data_vpu_req           ),
  .s_addr_a_i             ( data_vpu_addr          ),
  .s_be_a_i               ( data_vpu_be            ),
  .s_we_a_i               ( data_vpu_we            ),
  .s_wdata_a_i            ( data_vpu_wdata         ),

  .s_gnt_a_o              ( data_vpu_gnt           ),
  .s_rvalid_a_o           ( data_vpu_rvalid        ),
  .s_rdata_a_o            ( data_vpu_rdata         ),

  // input slave b cpu
  .s_req_b_i              ( data_cpu_req           ),
  .s_addr_b_i             ( data_cpu_addr          ),
  .s_be_b_i               ( data_cpu_be            ),
  .s_we_b_i               ( data_cpu_we            ),
  .s_wdata_b_i            ( data_cpu_wdata         ),

  .s_gnt_b_o              ( data_cpu_gnt           ),
  .s_rvalid_b_o           ( data_cpu_rvalid        ),
  .s_rdata_b_o            ( data_cpu_rdata         ),

  // output master
  .m_req_o                ( data_req              ),
  .m_addr_o               ( data_addr             ),
  .m_be_o                 ( data_be               ),
  .m_we_o                 ( data_we               ),
  .m_wdata_o              ( data_wdata            ),

  .m_gnt_i                ( data_gnt              ),
  .m_rvalid_i             ( data_rvalid           ),
  .m_rdata_i              ( data_rdata            )
);


// this handles read to RAM and memory mapped pseudo peripherals
mm_ram
#(.RAM_ADDR_WIDTH (RAM_ADDR_WIDTH),
  .INSTR_RDATA_WIDTH (INSTR_RDATA_WIDTH)
)
ram_i
(
  .clk_i          ( clk_i                          ),
  .rst_ni         ( rst_ni                         ),

  .instr_req_i    ( instr_req                      ),
  .instr_addr_i   ( instr_addr[RAM_ADDR_WIDTH-1:0] ),
  .instr_rdata_o  ( instr_rdata                    ),
  .instr_rvalid_o ( instr_rvalid                   ),
  .instr_gnt_o    ( instr_gnt                      ),

  .data_req_i     ( data_req                       ),
  .data_addr_i    ( data_addr                      ),
  .data_we_i      ( data_we                        ),
  .data_be_i      ( data_be                        ),
  .data_wdata_i   ( data_wdata                     ),
  .data_rdata_o   ( data_rdata                     ),
  .data_rvalid_o  ( data_rvalid                    ),
  .data_gnt_o     ( data_gnt                       ),

  .irq_id_i       ( irq_id_out                     ),
  .irq_ack_i      ( irq_ack                        ),
  .irq_id_o       ( irq_id_in                      ),
  .irq_o          ( irq                            ),

  .pc_core_id_i   ( riscv_core_i.pc_id             ),

  .tests_passed_o ( tests_passed_o                 ),
  .tests_failed_o ( tests_failed_o                 ),
  .exit_valid_o   ( exit_valid_o                   ),
  .exit_value_o   ( exit_value_o                   )
);

endmodule // riscv_wrapper
